module M (clk, data);
  input clk;
  output [31:0] data;
  reg [31:0] data;
endmodule
