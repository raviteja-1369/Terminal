module M (
  input wire clk,
  output reg [31:0] data
);
endmodule
